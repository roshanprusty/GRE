module filetest(in,out);
input [7:0] in;
output wire [7:0] out;
assign out = in;
endmodule