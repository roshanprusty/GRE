library verilog;
use verilog.vl_types.all;
entity t_ff_tb is
end t_ff_tb;
